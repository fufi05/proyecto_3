module module_decoabinbcd(
    input [7:0] b,
    output logic [7:0] bcd
);
always_comb begin
    case(b)
    // Binario sin signo a BCD
    8'b0000_0000: bcd = 8'b0000_0000; // 0
    8'b0000_0001: bcd = 8'b0000_0001; // 1
    8'b0000_0010: bcd = 8'b0000_0010; // 2
    8'b0000_0011: bcd = 8'b0000_0011; // 3
    8'b0000_0100: bcd = 8'b0000_0100; // 4
    8'b0000_0101: bcd = 8'b0000_0101; // 5
    8'b0000_0110: bcd = 8'b0000_0110; // 6
    8'b0000_0111: bcd = 8'b0000_0111; // 7
    8'b0000_1000: bcd = 8'b0000_1000; // 8
    8'b0000_1001: bcd = 8'b0000_1001; // 9
    8'b0000_1010: bcd = 8'b0001_0000; // 10
    8'b0000_1011: bcd = 8'b0001_0001; // 11
    8'b0000_1100: bcd = 8'b0001_0010; // 12
    8'b0000_1101: bcd = 8'b0001_0011; // 13
    8'b0000_1110: bcd = 8'b0001_0100; // 14
    8'b0000_1111: bcd = 8'b0001_0101; // 15
    8'b0001_0000: bcd = 8'b0001_0110; // 16
    8'b0001_0001: bcd = 8'b0001_0111; // 17
    8'b0001_0010: bcd = 8'b0001_1000; // 18
    8'b0001_0011: bcd = 8'b0001_1001; // 19
    8'b0001_0100: bcd = 8'b0010_0000; // 20
    8'b0001_0101: bcd = 8'b0010_0001; // 21
    8'b0001_0110: bcd = 8'b0010_0010; // 22
    8'b0001_0111: bcd = 8'b0010_0011; // 23
    8'b0001_1000: bcd = 8'b0010_0100; // 24
    8'b0001_1001: bcd = 8'b0010_0101; // 25
    8'b0001_1010: bcd = 8'b0010_0110; // 26
    8'b0001_1011: bcd = 8'b0010_0111; // 27
    8'b0001_1100: bcd = 8'b0010_1000; // 28
    8'b0001_1101: bcd = 8'b0010_1001; // 29
    8'b0001_1110: bcd = 8'b0011_0000; // 30
    8'b0001_1111: bcd = 8'b0011_0001; // 31
    8'b0010_0000: bcd = 8'b0011_0010; // 32
    8'b0010_0001: bcd = 8'b0011_0011; // 33
    8'b0010_0010: bcd = 8'b0011_0100; // 34
    8'b0010_0011: bcd = 8'b0011_0101; // 35
    8'b0010_0100: bcd = 8'b0011_0110; // 36
    8'b0010_0101: bcd = 8'b0011_0111; // 37
    8'b0010_0110: bcd = 8'b0011_1000; // 38
    8'b0010_0111: bcd = 8'b0011_1001; // 39
    8'b0010_1000: bcd = 8'b0100_0000; // 40
    8'b0010_1001: bcd = 8'b0100_0001; // 41
    8'b0010_1010: bcd = 8'b0100_0010; // 42
    8'b0010_1011: bcd = 8'b0100_0011; // 43
    8'b0010_1100: bcd = 8'b0100_0100; // 44
    8'b0010_1101: bcd = 8'b0100_0101; // 45
    8'b0010_1110: bcd = 8'b0100_0110; // 46
    8'b0010_1111: bcd = 8'b0100_0111; // 47
    8'b0011_0000: bcd = 8'b0100_1000; // 48
    8'b0011_0001: bcd = 8'b0100_1001; // 49
    8'b0011_0010: bcd = 8'b0101_0000; // 50
    8'b0011_0011: bcd = 8'b0101_0001; // 51
    8'b0011_0100: bcd = 8'b0101_0010; // 52
    8'b0011_0101: bcd = 8'b0101_0011; // 53
    8'b0011_0110: bcd = 8'b0101_0100; // 54
    8'b0011_0111: bcd = 8'b0101_0101; // 55
    8'b0011_1000: bcd = 8'b0101_0110; // 56
    8'b0011_1001: bcd = 8'b0101_0111; // 57
    8'b0011_1010: bcd = 8'b0101_1000; // 58
    8'b0011_1011: bcd = 8'b0101_1001; // 59
    8'b0011_1100: bcd = 8'b0110_0000; // 60
    8'b0011_1101: bcd = 8'b0110_0001; // 61
    8'b0011_1110: bcd = 8'b0110_0010; // 62
    8'b0011_1111: bcd = 8'b0110_0011; // 63
    8'b0100_0000: bcd = 8'b0110_0100; // 64
    8'b0100_0001: bcd = 8'b0110_0101; // 65
    8'b0100_0010: bcd = 8'b0110_0110; // 66
    8'b0100_0011: bcd = 8'b0110_0111; // 67
    8'b0100_0100: bcd = 8'b0110_1000; // 68
    8'b0100_0101: bcd = 8'b0110_1001; // 69
    8'b0100_0110: bcd = 8'b0111_0000; // 70
    8'b0100_0111: bcd = 8'b0111_0001; // 71
    8'b0100_1000: bcd = 8'b0111_0010; // 72
    8'b0100_1001: bcd = 8'b0111_0011; // 73
    8'b0100_1010: bcd = 8'b0111_0100; // 74
    8'b0100_1011: bcd = 8'b0111_0101; // 75
    8'b0100_1100: bcd = 8'b0111_0110; // 76
    8'b0100_1101: bcd = 8'b0111_0111; // 77
    8'b0100_1110: bcd = 8'b0111_1000; // 78
    8'b0100_1111: bcd = 8'b0111_1001; // 79
    8'b0101_0000: bcd = 8'b1000_0000; // 80
    8'b0101_0001: bcd = 8'b1000_0001; // 81
    default: bcd = 8'b00000000; // Default case to handle unexpected inputs
    endcase
end
endmodule