module module_multiplicador#(
    parameter N = 4
)(
    input logic clk,
    input logic rst,
    input logic [N-1:0] A,
    input logic [N-1:0] B,
    output logic [2*N-1:0] Y 
);

module_fsmbooth 
endmodule